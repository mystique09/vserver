module route