module middleware