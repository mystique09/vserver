module bootstrap

pub struct Env {}