module bootstrap

pub struct Database {}