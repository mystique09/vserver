module usecase