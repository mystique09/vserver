module repositories