module bootstrap

pub struct Application {}