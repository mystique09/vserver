module repository