module controller