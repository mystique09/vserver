module domain