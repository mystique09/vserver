module router